// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   cpu.u_reg_file
`define DMEM_PATH cpu.u_mem_control.u_dmem
`define IMEM_PATH cpu.u_mem_control.u_imem
`define BIOS_PATH cpu.u_mem_control.u_bios
`define CSR_PATH  cpu.u_mem_control.csr_reg
